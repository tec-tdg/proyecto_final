module MEMORYMAP(input logic  [6:0] dir,output logic [2:0] seleccion);
endmodule 
