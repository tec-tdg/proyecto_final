//Este procesador interpreta un ADD y  un ADD con inmediato

module CPU_V1();


endmodule