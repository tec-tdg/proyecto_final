module ADD_Instruction_TB();

endmodule